module shifter( dataA, dataB, Signal, dataOut );
input reset ;
input [31:0] dataA ;
input [31:0] dataB ; // sel
input [5:0] Signal ;
output [31:0] dataOut ;

wire[4:0] a ;
wire [31:0] temp ; // be the temp-result
wire[31:0] temp2 ;
wire[31:0] temp3 ;
wire[31:0] temp4 ;
wire[31:0] temp5 ;
wire[4:0] sel ;
assign a = dataB[4:0] ;
        
MUX2_1 mux01( .out( temp[0] ), .in0(1'b0) , .in1( dataA[0] ) , .sel(a[0] ) ) ;
MUX2_1 mux02( .out( temp[1] ), .in0(dataA[0]) , .in1( dataA[1] ) , .sel(a[0] ) ) ;
MUX2_1 mux03( .out( temp[2] ), .in0(dataA[1]) , .in1( dataA[2] ) , .sel(a[0] ) ) ;
MUX2_1 mux04( .out( temp[3] ), .in0(dataA[2]) , .in1( dataA[3] ) , .sel(a[0] ) ) ;
MUX2_1 mux05( .out( temp[4] ), .in0(dataA[3]) , .in1( dataA[4] ) , .sel(a[0] ) ) ;
MUX2_1 mux06( .out( temp[5] ), .in0(dataA[4]) , .in1( dataA[5] ) , .sel(a[0] ) ) ;
MUX2_1 mux07( .out( temp[6] ), .in0(dataA[5]) , .in1( dataA[6] ) , .sel(a[0] ) ) ;
MUX2_1 mux08( .out( temp[7] ), .in0(dataA[6]) , .in1( dataA[7] ) , .sel(a[0] ) ) ;
MUX2_1 mux09( .out( temp[8] ), .in0(dataA[7]) , .in1( dataA[8] ) , .sel(a[0] ) ) ;
MUX2_1 mux10( .out( temp[9] ), .in0(dataA[8]) , .in1( dataA[9] ) , .sel(a[0] ) ) ;
MUX2_1 mux11( .out( temp[10] ), .in0(dataA[9]) , .in1( dataA[10] ) , .sel(a[0] ) ) ;
MUX2_1 mux12( .out( temp[11] ), .in0(dataA[10]) , .in1( dataA[11] ) , .sel(a[0] ) ) ;
MUX2_1 mux13( .out( temp[12] ), .in0(dataA[11]) , .in1( dataA[12] ) , .sel(a[0] ) ) ;
MUX2_1 mux14( .out( temp[13] ), .in0(dataA[12]) , .in1( dataA[13] ) , .sel(a[0] ) ) ;
MUX2_1 mux15( .out( temp[14] ), .in0(dataA[13]) , .in1( dataA[14] ) , .sel(a[0] ) ) ;
MUX2_1 mux16( .out( temp[15] ), .in0(dataA[14]) , .in1( dataA[15] ) , .sel(a[0] ) ) ;
MUX2_1 mux17( .out( temp[16] ), .in0(dataA[15]) , .in1( dataA[16] ) , .sel(a[0] ) ) ;
MUX2_1 mux18( .out( temp[17] ), .in0(dataA[16]) , .in1( dataA[17] ) , .sel(a[0] ) ) ;
MUX2_1 mux19( .out( temp[18] ), .in0(dataA[17]) , .in1( dataA[18] ) , .sel(a[0] ) ) ;
MUX2_1 mux20( .out( temp[19] ), .in0(dataA[18]) , .in1( dataA[19] ) , .sel(a[0] ) ) ;
MUX2_1 mux21( .out( temp[20] ), .in0(dataA[19]) , .in1( dataA[20] ) , .sel(a[0] ) ) ;
MUX2_1 mux22( .out( temp[21] ), .in0(dataA[20]) , .in1( dataA[21] ) , .sel(a[0] ) ) ;
MUX2_1 mux23( .out( temp[22] ), .in0(dataA[21]) , .in1( dataA[22] ) , .sel(a[0] ) ) ;
MUX2_1 mux24( .out( temp[23] ), .in0(dataA[22]) , .in1( dataA[23] ) , .sel(a[0] ) ) ;
MUX2_1 mux25( .out( temp[24] ), .in0(dataA[23]) , .in1( dataA[24] ) , .sel(a[0] ) ) ;
MUX2_1 mux26( .out( temp[25] ), .in0(dataA[24]) , .in1( dataA[25] ) , .sel(a[0] ) ) ;
MUX2_1 mux27( .out( temp[26] ), .in0(dataA[25]) , .in1( dataA[26] ) , .sel(a[0] ) ) ;
MUX2_1 mux28( .out( temp[27] ), .in0(dataA[26]) , .in1( dataA[27] ) , .sel(a[0] ) ) ;
MUX2_1 mux29( .out( temp[28] ), .in0(dataA[27]) , .in1( dataA[28] ) , .sel(a[0] ) ) ;
MUX2_1 mux30( .out( temp[29] ), .in0(dataA[28]) , .in1( dataA[29] ) , .sel(a[0] ) ) ;
MUX2_1 mux31( .out( temp[30] ), .in0(dataA[29]) , .in1( dataA[30] ) , .sel(a[0] ) ) ;
MUX2_1 mux32( .out( temp[31] ), .in0(dataA[30]) , .in1( dataA[31] ) , .sel(a[0] ) ) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////
MUX2_1 mux001( .out( temp2[0] ), .in0(1'b0) , .in1( temp[0] ) , .sel(a[1] ) ) ;
MUX2_1 mux002( .out( temp2[1] ), .in0(1'b0) , .in1( temp[1] ) , .sel(a[1] ) ) ;
MUX2_1 mux003( .out( temp2[2] ), .in0(temp[0]) , .in1( temp[2] ) , .sel(a[1] ) ) ;
MUX2_1 mux004( .out( temp2[3] ), .in0(temp[1]) , .in1( temp[3] ) , .sel(a[1] ) ) ;
MUX2_1 mux005( .out( temp2[4] ), .in0(temp[2]) , .in1( temp[4] ) , .sel(a[1] ) ) ;
MUX2_1 mux006( .out( temp2[5] ), .in0(temp[3]) , .in1( temp[5] ) , .sel(a[1] ) ) ;
MUX2_1 mux007( .out( temp2[6] ), .in0(temp[4]) , .in1( temp[6] ) , .sel(a[1] ) ) ;
MUX2_1 mux008( .out( temp2[7] ), .in0(temp[5]) , .in1( temp[7] ) , .sel(a[1] ) ) ;
MUX2_1 mux009( .out( temp2[8] ), .in0(temp[6]) , .in1( temp[8] ) , .sel(a[1] ) ) ;
MUX2_1 mux010( .out( temp2[9] ), .in0(temp[7]) , .in1( temp[9] ) , .sel(a[1] ) ) ;
MUX2_1 mux011( .out( temp2[10] ), .in0(temp[8]) , .in1( temp[10] ) , .sel(a[1] ) ) ;
MUX2_1 mux012( .out( temp2[11] ), .in0(temp[9]) , .in1( temp[11] ) , .sel(a[1] ) ) ;
MUX2_1 mux013( .out( temp2[12] ), .in0(temp[10]) , .in1( temp[12] ) , .sel(a[1] ) ) ;
MUX2_1 mux014( .out( temp2[13] ), .in0(temp[11]) , .in1( temp[13] ) , .sel(a[1] ) ) ;
MUX2_1 mux015( .out( temp2[14] ), .in0(temp[12]) , .in1( temp[14] ) , .sel(a[1] ) ) ;
MUX2_1 mux016( .out( temp2[15] ), .in0(temp[13]) , .in1( temp[15] ) , .sel(a[1] ) ) ;
MUX2_1 mux017( .out( temp2[16] ), .in0(temp[14]) , .in1( temp[16] ) , .sel(a[1] ) ) ;
MUX2_1 mux018( .out( temp2[17] ), .in0(temp[15]) , .in1( temp[17] ) , .sel(a[1] ) ) ;
MUX2_1 mux019( .out( temp2[18] ), .in0(temp[16]) , .in1( temp[18] ) , .sel(a[1] ) ) ;
MUX2_1 mux020( .out( temp2[19] ), .in0(temp[17]) , .in1( temp[19] ) , .sel(a[1] ) ) ;
MUX2_1 mux021( .out( temp2[20] ), .in0(temp[18]) , .in1( temp[20] ) , .sel(a[1] ) ) ;
MUX2_1 mux022( .out( temp2[21] ), .in0(temp[19]) , .in1( temp[21] ) , .sel(a[1] ) ) ;
MUX2_1 mux023( .out( temp2[22] ), .in0(temp[20]) , .in1( temp[22] ) , .sel(a[1] ) ) ;
MUX2_1 mux024( .out( temp2[23] ), .in0(temp[21]) , .in1( temp[23] ) , .sel(a[1] ) ) ;
MUX2_1 mux025( .out( temp2[24] ), .in0(temp[22]) , .in1( temp[24] ) , .sel(a[1] ) ) ;
MUX2_1 mux026( .out( temp2[25] ), .in0(temp[23]) , .in1( temp[25] ) , .sel(a[1] ) ) ;
MUX2_1 mux027( .out( temp2[26] ), .in0(temp[24]) , .in1( temp[26] ) , .sel(a[1] ) ) ;
MUX2_1 mux028( .out( temp2[27] ), .in0(temp[25]) , .in1( temp[27] ) , .sel(a[1] ) ) ;
MUX2_1 mux029( .out( temp2[28] ), .in0(temp[26]) , .in1( temp[28] ) , .sel(a[1] ) ) ;
MUX2_1 mux030( .out( temp2[29] ), .in0(temp[27]) , .in1( temp[29] ) , .sel(a[1] ) ) ;
MUX2_1 mux031( .out( temp2[30] ), .in0(temp[28]) , .in1( temp[30] ) , .sel(a[1] ) ) ;
MUX2_1 mux032( .out( temp2[31] ), .in0(temp[29]) , .in1( temp[31] ) , .sel(a[1] ) ) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////
MUX2_1 mux0001( .out( temp3[0] ), .in0(1'b0) , .in1( temp2[0] ) , .sel(a[2] ) ) ;
MUX2_1 mux0002( .out( temp3[1] ), .in0(1'b0) , .in1( temp2[1] ) , .sel(a[2] ) ) ;
MUX2_1 mux0003( .out( temp3[2] ), .in0(1'b0) , .in1( temp2[2] ) , .sel(a[2] ) ) ;
MUX2_1 mux0004( .out( temp3[3] ), .in0(1'b0) , .in1( temp2[3] ) , .sel(a[2] ) ) ;
MUX2_1 mux0005( .out( temp3[4] ), .in0(temp2[0]) , .in1( temp2[4] ) , .sel(a[2] ) ) ;
MUX2_1 mux0006( .out( temp3[5] ), .in0(temp2[1]) , .in1( temp2[5] ) , .sel(a[2] ) ) ;
MUX2_1 mux0007( .out( temp3[6] ), .in0(temp2[2]) , .in1( temp2[6] ) , .sel(a[2] ) ) ;
MUX2_1 mux0008( .out( temp3[7] ), .in0(temp2[3]) , .in1( temp2[7] ) , .sel(a[2] ) ) ;
MUX2_1 mux0009( .out( temp3[8] ), .in0(temp2[4]) , .in1( temp2[8] ) , .sel(a[2] ) ) ;
MUX2_1 mux0010( .out( temp3[9] ), .in0(temp2[5]) , .in1( temp2[9] ) , .sel(a[2] ) ) ;
MUX2_1 mux0011( .out( temp3[10] ), .in0(temp2[6]) , .in1( temp2[10] ) , .sel(a[2] ) ) ;
MUX2_1 mux0012( .out( temp3[11] ), .in0(temp2[7]) , .in1( temp2[11] ) , .sel(a[2] ) ) ;
MUX2_1 mux0013( .out( temp3[12] ), .in0(temp2[8]) , .in1( temp2[12] ) , .sel(a[2] ) ) ;
MUX2_1 mux0014( .out( temp3[13] ), .in0(temp2[9]) , .in1( temp2[13] ) , .sel(a[2] ) ) ;
MUX2_1 mux0015( .out( temp3[14] ), .in0(temp2[10]) , .in1( temp2[14] ) , .sel(a[2] ) ) ;
MUX2_1 mux0016( .out( temp3[15] ), .in0(temp2[11]) , .in1( temp2[15] ) , .sel(a[2] ) ) ;
MUX2_1 mux0017( .out( temp3[16] ), .in0(temp2[12]) , .in1( temp2[16] ) , .sel(a[2] ) ) ;
MUX2_1 mux0018( .out( temp3[17] ), .in0(temp2[13]) , .in1( temp2[17] ) , .sel(a[2] ) ) ;
MUX2_1 mux0019( .out( temp3[18] ), .in0(temp2[14]) , .in1( temp2[18] ) , .sel(a[2] ) ) ;
MUX2_1 mux0020( .out( temp3[19] ), .in0(temp2[15]) , .in1( temp2[19] ) , .sel(a[2] ) ) ;
MUX2_1 mux0021( .out( temp3[20] ), .in0(temp2[16]) , .in1( temp2[20] ) , .sel(a[2] ) ) ;
MUX2_1 mux0022( .out( temp3[21] ), .in0(temp2[17]) , .in1( temp2[21] ) , .sel(a[2] ) ) ;
MUX2_1 mux0023( .out( temp3[22] ), .in0(temp2[18]) , .in1( temp2[22] ) , .sel(a[2] ) ) ;
MUX2_1 mux0024( .out( temp3[23] ), .in0(temp2[19]) , .in1( temp2[23] ) , .sel(a[2] ) ) ;
MUX2_1 mux0025( .out( temp3[24] ), .in0(temp2[20]) , .in1( temp2[24] ) , .sel(a[2] ) ) ;
MUX2_1 mux0026( .out( temp3[25] ), .in0(temp2[21]) , .in1( temp2[25] ) , .sel(a[2] ) ) ;
MUX2_1 mux0027( .out( temp3[26] ), .in0(temp2[22]) , .in1( temp2[26] ) , .sel(a[2] ) ) ;
MUX2_1 mux0028( .out( temp3[27] ), .in0(temp2[23]) , .in1( temp2[27] ) , .sel(a[2] ) ) ;
MUX2_1 mux0029( .out( temp3[28] ), .in0(temp2[24]) , .in1( temp2[28] ) , .sel(a[2] ) ) ;
MUX2_1 mux0030( .out( temp3[29] ), .in0(temp2[25]) , .in1( temp2[29] ) , .sel(a[2] ) ) ;
MUX2_1 mux0031( .out( temp3[30] ), .in0(temp2[26]) , .in1( temp2[30] ) , .sel(a[2] ) ) ;
MUX2_1 mux0032( .out( temp3[31] ), .in0(temp2[27]) , .in1( temp2[31] ) , .sel(a[2] ) ) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////
MUX2_1 mux00001( .out( temp4[0] ), .in0(1'b0) , .in1( temp3[0] ) , .sel(a[3] ) ) ;
MUX2_1 mux00002( .out( temp4[1] ), .in0(1'b0) , .in1( temp3[1] ) , .sel(a[3] ) ) ;
MUX2_1 mux00003( .out( temp4[2] ), .in0(1'b0) , .in1( temp3[2] ) , .sel(a[3] ) ) ;
MUX2_1 mux00004( .out( temp4[3] ), .in0(1'b0) , .in1( temp3[3] ) , .sel(a[3] ) ) ;
MUX2_1 mux00005( .out( temp4[4] ), .in0(1'b0) , .in1( temp3[4] ) , .sel(a[3] ) ) ;
MUX2_1 mux00006( .out( temp4[5] ), .in0(1'b0) , .in1( temp3[5] ) , .sel(a[3] ) ) ;
MUX2_1 mux00007( .out( temp4[6] ), .in0(1'b0) , .in1( temp3[6] ) , .sel(a[3] ) ) ;
MUX2_1 mux00008( .out( temp4[7] ), .in0(1'b0) , .in1( temp3[7] ) , .sel(a[3] ) ) ;
MUX2_1 mux00009( .out( temp4[8] ), .in0(temp3[0]) , .in1( temp3[8] ) , .sel(a[3] ) ) ;
MUX2_1 mux00010( .out( temp4[9] ), .in0(temp3[1]) , .in1( temp3[9] ) , .sel(a[3] ) ) ;
MUX2_1 mux00011( .out( temp4[10] ), .in0(temp3[2]) , .in1( temp3[10] ) , .sel(a[3] ) ) ;
MUX2_1 mux00012( .out( temp4[11] ), .in0(temp3[3]) , .in1( temp3[11] ) , .sel(a[3] ) ) ;
MUX2_1 mux00013( .out( temp4[12] ), .in0(temp3[4]) , .in1( temp3[12] ) , .sel(a[3] ) ) ;
MUX2_1 mux00014( .out( temp4[13] ), .in0(temp3[5]) , .in1( temp3[13] ) , .sel(a[3] ) ) ;
MUX2_1 mux00015( .out( temp4[14] ), .in0(temp3[6]) , .in1( temp3[14] ) , .sel(a[3] ) ) ;
MUX2_1 mux00016( .out( temp4[15] ), .in0(temp3[7]) , .in1( temp3[15] ) , .sel(a[3] ) ) ;
MUX2_1 mux00017( .out( temp4[16] ), .in0(temp3[8]) , .in1( temp3[16] ) , .sel(a[3] ) ) ;
MUX2_1 mux00018( .out( temp4[17] ), .in0(temp3[9]) , .in1( temp3[17] ) , .sel(a[3] ) ) ;
MUX2_1 mux00019( .out( temp4[18] ), .in0(temp3[10]) , .in1( temp3[18] ) , .sel(a[3] ) ) ;
MUX2_1 mux00020( .out( temp4[19] ), .in0(temp3[11]) , .in1( temp3[19] ) , .sel(a[3] ) ) ;
MUX2_1 mux00021( .out( temp4[20] ), .in0(temp3[12]) , .in1( temp3[20] ) , .sel(a[3] ) ) ;
MUX2_1 mux00022( .out( temp4[21] ), .in0(temp3[13]) , .in1( temp3[21] ) , .sel(a[3] ) ) ;
MUX2_1 mux00023( .out( temp4[22] ), .in0(temp3[14]) , .in1( temp3[22] ) , .sel(a[3] ) ) ;
MUX2_1 mux00024( .out( temp4[23] ), .in0(temp3[15]) , .in1( temp3[23] ) , .sel(a[3] ) ) ;
MUX2_1 mux00025( .out( temp4[24] ), .in0(temp3[16]) , .in1( temp3[24] ) , .sel(a[3] ) ) ;
MUX2_1 mux00026( .out( temp4[25] ), .in0(temp3[17]) , .in1( temp3[25] ) , .sel(a[3] ) ) ;
MUX2_1 mux00027( .out( temp4[26] ), .in0(temp3[18]) , .in1( temp3[26] ) , .sel(a[3] ) ) ;
MUX2_1 mux00028( .out( temp4[27] ), .in0(temp3[19]) , .in1( temp3[27] ) , .sel(a[3] ) ) ;
MUX2_1 mux00029( .out( temp4[28] ), .in0(temp3[20]) , .in1( temp3[28] ) , .sel(a[3] ) ) ;
MUX2_1 mux00030( .out( temp4[29] ), .in0(temp3[21]) , .in1( temp3[29] ) , .sel(a[3] ) ) ;
MUX2_1 mux00031( .out( temp4[30] ), .in0(temp3[22]) , .in1( temp3[30] ) , .sel(a[3] ) ) ;
MUX2_1 mux00032( .out( temp4[31] ), .in0(temp3[23]) , .in1( temp3[31] ) , .sel(a[3] ) ) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////
MUX2_1 mux000001( .out( temp5[0] ), .in0(1'b0) , .in1( temp4[0] ) , .sel(a[4] ) ) ;
MUX2_1 mux000002( .out( temp5[1] ), .in0(1'b0) , .in1( temp4[1] ) , .sel(a[4] ) ) ;
MUX2_1 mux000003( .out( temp5[2] ), .in0(1'b0) , .in1( temp4[2] ) , .sel(a[4] ) ) ;
MUX2_1 mux000004( .out( temp5[3] ), .in0(1'b0) , .in1( temp4[3] ) , .sel(a[4] ) ) ;
MUX2_1 mux000005( .out( temp5[4] ), .in0(1'b0) , .in1( temp4[4] ) , .sel(a[4] ) ) ;
MUX2_1 mux000006( .out( temp5[5] ), .in0(1'b0) , .in1( temp4[5] ) , .sel(a[4] ) ) ;
MUX2_1 mux000007( .out( temp5[6] ), .in0(1'b0) , .in1( temp4[6] ) , .sel(a[4] ) ) ;
MUX2_1 mux000008( .out( temp5[7] ), .in0(1'b0) , .in1( temp4[7] ) , .sel(a[4] ) ) ;
MUX2_1 mux000009( .out( temp5[8] ), .in0(1'b0) , .in1( temp4[8] ) , .sel(a[4] ) ) ;
MUX2_1 mux000010( .out( temp5[9] ), .in0(1'b0) , .in1( temp4[9] ) , .sel(a[4] ) ) ;
MUX2_1 mux000011( .out( temp5[10] ), .in0(1'b0) , .in1( temp4[10] ) , .sel(a[4] ) ) ;
MUX2_1 mux000012( .out( temp5[11] ), .in0(1'b0) , .in1( temp4[11] ) , .sel(a[4] ) ) ;
MUX2_1 mux000013( .out( temp5[12] ), .in0(1'b0) , .in1( temp4[12] ) , .sel(a[4] ) ) ;
MUX2_1 mux000014( .out( temp5[13] ), .in0(1'b0) , .in1( temp4[13] ) , .sel(a[4] ) ) ;
MUX2_1 mux000015( .out( temp5[14] ), .in0(1'b0) , .in1( temp4[14] ) , .sel(a[4] ) ) ;
MUX2_1 mux000016( .out( temp5[15] ), .in0(1'b0) , .in1( temp4[15] ) , .sel(a[4] ) ) ;
MUX2_1 mux000017( .out( temp5[16] ), .in0(temp4[0]) , .in1( temp4[16] ) , .sel(a[4] ) ) ;
MUX2_1 mux000018( .out( temp5[17] ), .in0(temp4[1]) , .in1( temp4[17] ) , .sel(a[4] ) ) ;
MUX2_1 mux000019( .out( temp5[18] ), .in0(temp4[2]) , .in1( temp4[18] ) , .sel(a[4] ) ) ;
MUX2_1 mux000020( .out( temp5[19] ), .in0(temp4[4]) , .in1( temp4[19] ) , .sel(a[4] ) ) ;
MUX2_1 mux000021( .out( temp5[20] ), .in0(temp4[4]) , .in1( temp4[20] ) , .sel(a[4] ) ) ;
MUX2_1 mux000022( .out( temp5[21] ), .in0(temp4[5]) , .in1( temp4[21] ) , .sel(a[4] ) ) ;
MUX2_1 mux000023( .out( temp5[22] ), .in0(temp4[6]) , .in1( temp4[22] ) , .sel(a[4] ) ) ;
MUX2_1 mux000024( .out( temp5[23] ), .in0(temp4[7]) , .in1( temp4[23] ) , .sel(a[4] ) ) ;
MUX2_1 mux000025( .out( temp5[24] ), .in0(temp4[8]) , .in1( temp4[24] ) , .sel(a[4] ) ) ;
MUX2_1 mux000026( .out( temp5[25] ), .in0(temp4[9]) , .in1( temp4[25] ) , .sel(a[4] ) ) ;
MUX2_1 mux000027( .out( temp5[26] ), .in0(temp4[10]) , .in1( temp4[26] ) , .sel(a[4] ) ) ;
MUX2_1 mux000028( .out( temp5[27] ), .in0(temp4[11]) , .in1( temp4[27] ) , .sel(a[4] ) ) ;
MUX2_1 mux000029( .out( temp5[28] ), .in0(temp4[12]) , .in1( temp4[28] ) , .sel(a[4] ) ) ;
MUX2_1 mux000030( .out( temp5[29] ), .in0(temp4[13]) , .in1( temp4[29] ) , .sel(a[4] ) ) ;
MUX2_1 mux000031( .out( temp5[30] ), .in0(temp4[14]) , .in1( temp4[30] ) , .sel(a[4] ) ) ;
MUX2_1 mux000032( .out( temp5[31] ), .in0(temp4[15]) , .in1( temp4[31] ) , .sel(a[4] ) ) ;
/////////////////////////////////////////////////////////////////////////////////////////////////////////
assign dataOut = temp5 ;

endmodule